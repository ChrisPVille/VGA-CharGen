//640x480@60Hz definitions (80 col text)

parameter H_ACTIVE = 640;
parameter H_FP = 16;
parameter H_SYN = 96;
parameter H_BP = 48;
parameter V_ACTIVE = 480;
parameter V_FP = 10;
parameter V_SYN = 2;
parameter V_BP = 29;

parameter N_COL = 80;
parameter N_ROW = 30;