//1920x1080@60Hz definitions (240 col text)

parameter H_ACTIVE = 1920;
parameter H_FP = 88;
parameter H_SYN = 44;
parameter H_BP = 148;
parameter V_ACTIVE = 1080;
parameter V_FP = 4;
parameter V_SYN = 5;
parameter V_BP = 36;

parameter N_COL = 240;
parameter N_ROW = 68;